.title KiCad schematic
.include "models/BZX84C4V7.spice.txt"
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/CGJ4C2C0G2A101J060AA_p.mod"
.include "models/ZXCT1082.spice.txt"
XU4 /COCM 0 /SP /SN VDD ZXCT1082
XU5 /SP /SN CGJ4C2C0G2A101J060AA_p
R4 /SN /PWR_OUT 2.74k
R5 /PWR_IN /PWR_OUT 0.1
R6 /PWR_IN /PWR_OUT 0.1
R3 /SP /PWR_IN 2.74k
I1 /PWR_OUT 0 {ILOAD}
V2 /PWR_IN 0 {VSOURCE}
R2 /COCM 0 68.1k
V1 VDD 0 {VSUPPLY}
R1 /OUT /COCM 100
XU2 /OUT 0 C2012C0G2A102J060AA_p
XU1 0 /OUT DI_BZX84C4V7
XU3 VDD 0 C2012X7R2A104K125AA_p
.end
